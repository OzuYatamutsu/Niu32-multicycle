module RegisterFile(regOutput);
    reg [(DBITS - 1):0] regs[31:0];
    
endmodule

