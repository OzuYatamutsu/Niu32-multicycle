library verilog;
use verilog.vl_types.all;
entity Niu32_multicycle is
    generic(
        WORD_SIZE       : integer := 32;
        INSTR_SIZE      : integer := 4;
        IMM_SIZE        : integer := 17;
        NUM_REGS        : integer := 32;
        REG_BITS        : integer := 5;
        OP_BITS         : integer := 5;
        STATE_BITS      : integer := 6;
        ADDR_HEX        : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_LEDR       : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_LEDG       : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_KEY        : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_SWITCH     : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_MIF        : string  := "test1.mif";
        IMEM_WORDS      : integer := 2048;
        DMEM_WORDS      : integer := 2048;
        MEM_ADDR_BITS   : integer := 13;
        MEM_WORD_OFFSET : integer := 2;
        PC_STARTLOC     : integer := 0;
        BUS_NOSIG       : vl_notype;
        BYTE_SEL_MASK   : vl_notype;
        OP1_ALUI        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        OP1_ADDI        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        OP1_MLTI        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        OP1_DIVI        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        OP1_ANDI        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        OP1_ORI         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        OP1_XORI        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        OP1_SULI        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        OP1_SSLI        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        OP1_SURI        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        OP1_SSRI        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        OP1_LW          : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        OP1_LB          : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        OP1_SW          : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi1);
        OP1_SB          : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi0);
        OP1_LUI         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi0);
        OP1_BEQ         : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi0, Hi0);
        OP1_BNE         : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi0, Hi1);
        OP1_BLT         : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi1, Hi0);
        OP1_BLE         : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi1, Hi1);
        OP1_JAL         : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi1);
        OP2_SUB         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        OP2_ADD         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        OP2_MLT         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        OP2_DIV         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        OP2_NOT         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        OP2_AND         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        OP2_OR          : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        OP2_XOR         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        OP2_SUL         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        OP2_SSL         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        OP2_SUR         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        OP2_SSR         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        OP2_EQ          : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        OP2_NEQ         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        OP2_LT          : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi0);
        OP2_LEQ         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi1);
        OP3_LUI         : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi0, Hi0);
        OP3_BITSEL      : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi0, Hi1);
        OP3_BITUNSET    : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi0);
        OP3_BITSET      : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi1);
        S_FETCH         : vl_logic_vector;
        S_DECODE        : vl_logic_vector;
        S_ALU0I         : vl_logic_vector;
        S_ALU0R         : vl_logic_vector;
        S_ALU1          : vl_logic_vector;
        S_ALU2          : vl_logic_vector;
        S_ALU3          : vl_logic_vector;
        S_LW0           : vl_logic_vector;
        S_LW1           : vl_logic_vector;
        S_LW2           : vl_logic_vector;
        S_LW3           : vl_logic_vector;
        S_LB0           : vl_logic_vector;
        S_LB1           : vl_logic_vector;
        S_LB2           : vl_logic_vector;
        S_LB3           : vl_logic_vector;
        S_SW0           : vl_logic_vector;
        S_SW1           : vl_logic_vector;
        S_SW2           : vl_logic_vector;
        S_SW3           : vl_logic_vector;
        S_SB0           : vl_logic_vector;
        S_SB1           : vl_logic_vector;
        S_SB2           : vl_logic_vector;
        S_SB3           : vl_logic_vector;
        S_SB4           : vl_logic_vector;
        S_SB5           : vl_logic_vector;
        S_LUI0          : vl_logic_vector;
        S_LUI1          : vl_logic_vector;
        S_LUI2          : vl_logic_vector;
        S_BRCH0         : vl_logic_vector;
        S_BRCH1         : vl_logic_vector;
        S_BRCH2         : vl_logic_vector;
        S_BRCH3         : vl_logic_vector;
        S_BRCH4         : vl_logic_vector;
        S_BRCH5         : vl_logic_vector;
        S_JUMP0         : vl_logic_vector;
        S_JUMP1         : vl_logic_vector;
        S_ERROR         : vl_logic_vector;
        \ON\            : vl_logic := Hi1;
        OFF             : vl_logic := Hi0
    );
    port(
        SWITCH          : in     vl_logic_vector(9 downto 0);
        KEY             : in     vl_logic_vector(3 downto 0);
        LEDR            : out    vl_logic_vector(9 downto 0);
        LEDG            : out    vl_logic_vector(7 downto 0);
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        CLOCK_50        : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of WORD_SIZE : constant is 1;
    attribute mti_svvh_generic_type of INSTR_SIZE : constant is 1;
    attribute mti_svvh_generic_type of IMM_SIZE : constant is 1;
    attribute mti_svvh_generic_type of NUM_REGS : constant is 1;
    attribute mti_svvh_generic_type of REG_BITS : constant is 1;
    attribute mti_svvh_generic_type of OP_BITS : constant is 1;
    attribute mti_svvh_generic_type of STATE_BITS : constant is 1;
    attribute mti_svvh_generic_type of ADDR_HEX : constant is 1;
    attribute mti_svvh_generic_type of ADDR_LEDR : constant is 1;
    attribute mti_svvh_generic_type of ADDR_LEDG : constant is 1;
    attribute mti_svvh_generic_type of ADDR_KEY : constant is 1;
    attribute mti_svvh_generic_type of ADDR_SWITCH : constant is 1;
    attribute mti_svvh_generic_type of INIT_MIF : constant is 1;
    attribute mti_svvh_generic_type of IMEM_WORDS : constant is 1;
    attribute mti_svvh_generic_type of DMEM_WORDS : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADDR_BITS : constant is 1;
    attribute mti_svvh_generic_type of MEM_WORD_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PC_STARTLOC : constant is 1;
    attribute mti_svvh_generic_type of BUS_NOSIG : constant is 3;
    attribute mti_svvh_generic_type of BYTE_SEL_MASK : constant is 3;
    attribute mti_svvh_generic_type of OP1_ALUI : constant is 1;
    attribute mti_svvh_generic_type of OP1_ADDI : constant is 1;
    attribute mti_svvh_generic_type of OP1_MLTI : constant is 1;
    attribute mti_svvh_generic_type of OP1_DIVI : constant is 1;
    attribute mti_svvh_generic_type of OP1_ANDI : constant is 1;
    attribute mti_svvh_generic_type of OP1_ORI : constant is 1;
    attribute mti_svvh_generic_type of OP1_XORI : constant is 1;
    attribute mti_svvh_generic_type of OP1_SULI : constant is 1;
    attribute mti_svvh_generic_type of OP1_SSLI : constant is 1;
    attribute mti_svvh_generic_type of OP1_SURI : constant is 1;
    attribute mti_svvh_generic_type of OP1_SSRI : constant is 1;
    attribute mti_svvh_generic_type of OP1_LW : constant is 1;
    attribute mti_svvh_generic_type of OP1_LB : constant is 1;
    attribute mti_svvh_generic_type of OP1_SW : constant is 1;
    attribute mti_svvh_generic_type of OP1_SB : constant is 1;
    attribute mti_svvh_generic_type of OP1_LUI : constant is 1;
    attribute mti_svvh_generic_type of OP1_BEQ : constant is 1;
    attribute mti_svvh_generic_type of OP1_BNE : constant is 1;
    attribute mti_svvh_generic_type of OP1_BLT : constant is 1;
    attribute mti_svvh_generic_type of OP1_BLE : constant is 1;
    attribute mti_svvh_generic_type of OP1_JAL : constant is 1;
    attribute mti_svvh_generic_type of OP2_SUB : constant is 1;
    attribute mti_svvh_generic_type of OP2_ADD : constant is 1;
    attribute mti_svvh_generic_type of OP2_MLT : constant is 1;
    attribute mti_svvh_generic_type of OP2_DIV : constant is 1;
    attribute mti_svvh_generic_type of OP2_NOT : constant is 1;
    attribute mti_svvh_generic_type of OP2_AND : constant is 1;
    attribute mti_svvh_generic_type of OP2_OR : constant is 1;
    attribute mti_svvh_generic_type of OP2_XOR : constant is 1;
    attribute mti_svvh_generic_type of OP2_SUL : constant is 1;
    attribute mti_svvh_generic_type of OP2_SSL : constant is 1;
    attribute mti_svvh_generic_type of OP2_SUR : constant is 1;
    attribute mti_svvh_generic_type of OP2_SSR : constant is 1;
    attribute mti_svvh_generic_type of OP2_EQ : constant is 1;
    attribute mti_svvh_generic_type of OP2_NEQ : constant is 1;
    attribute mti_svvh_generic_type of OP2_LT : constant is 1;
    attribute mti_svvh_generic_type of OP2_LEQ : constant is 1;
    attribute mti_svvh_generic_type of OP3_LUI : constant is 1;
    attribute mti_svvh_generic_type of OP3_BITSEL : constant is 1;
    attribute mti_svvh_generic_type of OP3_BITUNSET : constant is 1;
    attribute mti_svvh_generic_type of OP3_BITSET : constant is 1;
    attribute mti_svvh_generic_type of S_FETCH : constant is 4;
    attribute mti_svvh_generic_type of S_DECODE : constant is 4;
    attribute mti_svvh_generic_type of S_ALU0I : constant is 4;
    attribute mti_svvh_generic_type of S_ALU0R : constant is 4;
    attribute mti_svvh_generic_type of S_ALU1 : constant is 4;
    attribute mti_svvh_generic_type of S_ALU2 : constant is 4;
    attribute mti_svvh_generic_type of S_ALU3 : constant is 4;
    attribute mti_svvh_generic_type of S_LW0 : constant is 4;
    attribute mti_svvh_generic_type of S_LW1 : constant is 4;
    attribute mti_svvh_generic_type of S_LW2 : constant is 4;
    attribute mti_svvh_generic_type of S_LW3 : constant is 4;
    attribute mti_svvh_generic_type of S_LB0 : constant is 4;
    attribute mti_svvh_generic_type of S_LB1 : constant is 4;
    attribute mti_svvh_generic_type of S_LB2 : constant is 4;
    attribute mti_svvh_generic_type of S_LB3 : constant is 4;
    attribute mti_svvh_generic_type of S_SW0 : constant is 4;
    attribute mti_svvh_generic_type of S_SW1 : constant is 4;
    attribute mti_svvh_generic_type of S_SW2 : constant is 4;
    attribute mti_svvh_generic_type of S_SW3 : constant is 4;
    attribute mti_svvh_generic_type of S_SB0 : constant is 4;
    attribute mti_svvh_generic_type of S_SB1 : constant is 4;
    attribute mti_svvh_generic_type of S_SB2 : constant is 4;
    attribute mti_svvh_generic_type of S_SB3 : constant is 4;
    attribute mti_svvh_generic_type of S_SB4 : constant is 4;
    attribute mti_svvh_generic_type of S_SB5 : constant is 4;
    attribute mti_svvh_generic_type of S_LUI0 : constant is 4;
    attribute mti_svvh_generic_type of S_LUI1 : constant is 4;
    attribute mti_svvh_generic_type of S_LUI2 : constant is 4;
    attribute mti_svvh_generic_type of S_BRCH0 : constant is 4;
    attribute mti_svvh_generic_type of S_BRCH1 : constant is 4;
    attribute mti_svvh_generic_type of S_BRCH2 : constant is 4;
    attribute mti_svvh_generic_type of S_BRCH3 : constant is 4;
    attribute mti_svvh_generic_type of S_BRCH4 : constant is 4;
    attribute mti_svvh_generic_type of S_BRCH5 : constant is 4;
    attribute mti_svvh_generic_type of S_JUMP0 : constant is 4;
    attribute mti_svvh_generic_type of S_JUMP1 : constant is 4;
    attribute mti_svvh_generic_type of S_ERROR : constant is 4;
    attribute mti_svvh_generic_type of \ON\ : constant is 1;
    attribute mti_svvh_generic_type of OFF : constant is 1;
end Niu32_multicycle;
